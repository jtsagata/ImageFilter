LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE constants IS
	CONSTANT MSIZE : NATURAL := 4;
	-- 4 bit X 8 bit + sign
	CONSTANT MRESULT : NATURAL := 13;
END constants;

PACKAGE BODY constants IS

END constants;
